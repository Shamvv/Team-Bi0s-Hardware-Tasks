* example.sch
* DSCH 2.7a
* created 16-04-2022 10.36.34 AM
*
* Input button "in1" 2
VBTN1 2 0 DC 0 PULSE(0 1.2 1.00N 0.1N 0.1N 1.00N 3.00N )
* Output "out1" 16
* Input button "in2" 4
VBTN2 4 0 DC 0 PULSE(0 1.2 2.00N 0.1N 0.1N 2.00N 5.00N )
* Input button "in3" 6
VBTN3 6 0 DC 0 PULSE(0 1.2 3.00N 0.1N 0.1N 3.00N 7.00N )
* Input button "in4" 8
VBTN4 8 0 DC 0 PULSE(0 1.2 4.00N 0.1N 0.1N 4.00N 9.00N )
*
* Mos models in 0.12µm
* Model 3 n-channel MOS
.MODEL  TN  NMOS
+ LEVEL=3            TPG=+1
+ GAMMA=0.2          THETA=0.5          KAPPA=0.1        ETA=0.002
+ DELTA=0.0          UO=620             VMAX=100E3       VTO=0.35
+ TOX=3e-9           XJ=0.1U            LD=0.00U         NSUB=1E+18
+ NSS=0.2            NFS=7E11
+ CJ=4.091E-4        MJ=0.307           PB=1.0
+ CJSW=3.078E-10     MJSW=1.0E-2
+ CGSO=3.93E-10      CGDO=3.93E-10
* Model 3 p-channel MOS
.MODEL  TP  PMOS
+ LEVEL=3            TPG=-1
+ GAMMA=0.2          THETA=0.5          KAPPA=0.01         ETA=0.001
+ DELTA=0.0          UO=250             VMAX=500E3         VTO=-0.35
+ TOX=3E-9          XJ=0.1U             LD=0.0U             NSUB=1E+18
+ NSS=0.0            NFS=7E11
+ CJ=6.852E-4        MJ=0.429           PB=1.0
+ CJSW=5.217E-10     MJSW=0.351
+ CGSO=7.29E-10      CGDO=7.29E-10
.TRAN 0.1N 50N
* Commands for WinSpice3
* No break in output file
*#set nobreak
* Dump time and volts in "out.txt"
*#print V(2) V(4) V(6) V(8)  V(16)  > out.txt
* Run simulation
*#run
* Show the result in a window
*#plot V(2) V(4) V(6) V(8)  V(16) 
.OPTIONS DELMIN=0 RELTOL=1E-6
.END
